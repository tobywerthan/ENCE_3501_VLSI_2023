*** SPICE deck for cell buftri_c_1x_sim{lay} from library Werthan_ALU
*** Created on Mon Nov 13, 2023 00:13:23
*** Last revised on Tue Nov 14, 2023 15:39:07
*** Written on Tue Nov 14, 2023 15:40:20 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_ALU__buftri_c_1x FROM CELL buftri_c_1x{lay}
.SUBCKT Werthan_ALU__buftri_c_1x d en gnd vdd y
Mnmos@0 net@62 en gnd gnd N_1u L=0.6U W=1.8U AS=6.54P AD=3.375P PS=17.4U PD=7.5U
Mnmos@2 net@73 en y gnd N_1u L=0.6U W=4.2U AS=7.65P AD=2.228P PS=13.2U PD=5.85U
Mnmos@3 gnd net@119 net@73 gnd N_1u L=0.6U W=4.2U AS=2.228P AD=6.54P PS=5.85U PD=17.4U
Mnmos@6 net@119 d gnd gnd N_1u L=0.6U W=1.8U AS=6.54P AD=3.375P PS=17.4U PD=7.5U
Mpmos@0 net@62 en vdd vdd P_1u L=0.6U W=2.7U AS=7.98P AD=3.375P PS=19.2U PD=7.5U
Mpmos@2 net@64 net@62 y vdd P_1u L=0.6U W=6U AS=7.65P AD=3.038P PS=13.2U PD=7.65U
Mpmos@3 vdd net@119 net@64 vdd P_1u L=0.6U W=6U AS=3.038P AD=7.98P PS=7.65U PD=19.2U
Mpmos@5 net@119 d vdd vdd P_1u L=0.6U W=2.7U AS=7.98P AD=3.375P PS=19.2U PD=7.5U
.ENDS Werthan_ALU__buftri_c_1x

*** TOP LEVEL CELL: buftri_c_1x_sim{lay}
Xbuftri_c@0 d en gnd vdd y Werthan_ALU__buftri_c_1x

* Spice Code nodes in cell cell 'buftri_c_1x_sim{lay}'
vdd vdd 0 dc 5
ven en 0 dc 5
vd d 0 pulse(0v 5v 0 1n 1n 10n 20n) 
.tran 0 60n
.include cmosedu_models.txt
.END

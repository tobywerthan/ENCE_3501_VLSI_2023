*** SPICE deck for cell charge_pump_3_stage_sim{sch} from library Werthan_DC_to_DC
*** Created on Wed Nov 08, 2023 21:44:42
*** Last revised on Sat Nov 11, 2023 19:16:24
*** Written on Sat Nov 11, 2023 19:30:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_DC_to_DC__charge_pump_3_stage FROM CELL charge_pump_3_stage{sch}
.SUBCKT Werthan_DC_to_DC__charge_pump_3_stage osc osc2 vout
** GLOBAL gnd
** GLOBAL vdd
Ccap@0 osc net@136 100u
Ccap@1 osc2 net@133 100u
Ccap@2 osc net@130 100u
Ccap@3 gnd vout 100u
Mnmos@0 vdd vdd net@136 gnd N_50n L=0.3U W=3U
Mnmos@1 net@136 net@136 net@133 gnd N_50n L=0.3U W=3U
Mnmos@2 net@133 net@133 net@130 gnd N_50n L=0.3U W=3U
Mnmos@3 net@130 net@130 vout gnd N_50n L=0.3U W=3U
Rresnwell@0 vout gnd 2MEG
.ENDS Werthan_DC_to_DC__charge_pump_3_stage

.global gnd vdd

*** TOP LEVEL CELL: charge_pump_3_stage_sim{sch}
Xcharge_p@0 osc osc2 vout Werthan_DC_to_DC__charge_pump_3_stage

* Spice Code nodes in cell cell 'charge_pump_3_stage_sim{sch}'
vdd vdd 0 DC 1v
vosc osc 0 pulse(0v 1v 0 1p 1p 0.025 0.05)
vosc2 osc2 0 pulse(0v 1v 0.025 1p 1p 0.025 0.05)
.tran 0 1000 1m
.include cmosedu_models.txt
.END

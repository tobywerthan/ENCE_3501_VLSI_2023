*** SPICE deck for cell ring_oscillator{sch} from library Werthan_DC_to_DC
*** Created on Thu Nov 09, 2023 15:32:22
*** Last revised on Sat Nov 11, 2023 10:39:42
*** Written on Sat Nov 11, 2023 10:39:56 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_DC_to_DC__NAND FROM CELL Werthan_DC_to_DC:NAND{sch}
.SUBCKT Werthan_DC_to_DC__NAND A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A net@11 gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@11 B gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 Y A vdd vdd PMOS L=0.6U W=1.8U
Mpmos@2 Y B vdd vdd PMOS L=0.6U W=1.8U
.ENDS Werthan_DC_to_DC__NAND

*** SUBCIRCUIT Werthan_DC_to_DC__NOT FROM CELL Werthan_DC_to_DC:NOT{sch}
.SUBCKT Werthan_DC_to_DC__NOT A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 Y A vdd vdd PMOS L=0.6U W=1.8U
.ENDS Werthan_DC_to_DC__NOT

.global gnd vdd

*** TOP LEVEL CELL: Werthan_DC_to_DC:ring_oscillator{sch}
Ccap@0 gnd net@59 10u
Ccap@1 gnd net@65 10u
Ccap@2 gnd net@71 10u
XNAND@0 En osc net@59 Werthan_DC_to_DC__NAND
XNOT@0 net@59 net@71 Werthan_DC_to_DC__NOT
XNOT@1 net@71 net@65 Werthan_DC_to_DC__NOT
XNOT@2 net@65 osc2 Werthan_DC_to_DC__NOT
XNOT@3 osc2 osc Werthan_DC_to_DC__NOT

* Spice Code nodes in cell cell 'Werthan_DC_to_DC:ring_oscillator{sch}'
vdd vdd 0 DC 5v
vin d_in 0 pulse(0v 5v 10n 1n 1n 40n 40n)
.tran 0 40n
.include cmosedu_models.txt
.END

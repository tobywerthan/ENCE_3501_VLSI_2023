*** SPICE deck for cell NAND_sim{sch} from library Werthan_full_adder
*** Created on Fri Oct 20, 2023 10:05:23
*** Last revised on Fri Oct 27, 2023 11:41:59
*** Written on Fri Oct 27, 2023 11:42:02 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_full_adder__NAND FROM CELL NAND{sch}
.SUBCKT Werthan_full_adder__NAND A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A net@11 gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@11 B gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 Y A vdd vdd PMOS L=0.6U W=1.8U
Mpmos@2 Y B vdd vdd PMOS L=0.6U W=1.8U
.ENDS Werthan_full_adder__NAND

.global gnd vdd

*** TOP LEVEL CELL: NAND_sim{sch}
XNAND@0 in vdd out Werthan_full_adder__NAND

* Spice Code nodes in cell cell 'NAND_sim{sch}'
vdd vdd 0 DC 5
vin in 0 pulse(0v 5v 10n 1n 1n 40n 40n)
.tran 0 40n
.include C5_models.txt
.END

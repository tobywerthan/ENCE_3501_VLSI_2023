*** SPICE deck for cell ring_oscillator_sim{sch} from library Werthan_Ring_Oscillator
*** Created on Wed Nov 01, 2023 11:48:57
*** Last revised on Wed Nov 01, 2023 11:49:54
*** Written on Wed Nov 08, 2023 21:47:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_Ring_Oscillator__NOT_gate FROM CELL NOT_gate{sch}
.SUBCKT Werthan_Ring_Oscillator__NOT_gate A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd N_1u L=0.6U W=3U
Mpmos@0 Y A vdd vdd P_1u L=0.6U W=6U
.ENDS Werthan_Ring_Oscillator__NOT_gate

*** SUBCIRCUIT Werthan_Ring_Oscillator__ring_oscillator FROM CELL ring_oscillator{sch}
.SUBCKT Werthan_Ring_Oscillator__ring_oscillator osc_out
** GLOBAL gnd
** GLOBAL vdd
XNOT_gate@0 osc_out net@0 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@1 net@0 net@1 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@2 net@1 net@2 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@3 net@2 net@6 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@11 net@6 net@3 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@12 net@3 net@4 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@13 net@4 net@5 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@14 net@5 net@9 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@15 net@9 net@7 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@16 net@7 net@8 Werthan_Ring_Oscillator__NOT_gate
XNOT_gate@17 net@8 osc_out Werthan_Ring_Oscillator__NOT_gate
.ENDS Werthan_Ring_Oscillator__ring_oscillator

.global gnd vdd

*** TOP LEVEL CELL: ring_oscillator_sim{sch}
Xring_osc@0 osc_out Werthan_Ring_Oscillator__ring_oscillator

* Spice Code nodes in cell cell 'ring_oscillator_sim{sch}'
vdd vdd 0 DC 5v
vin d_in 0 pulse(0v 5v 10n 1n 1n 40n 40n)
.tran 0 40n
.include cmosedu_models.txt
.END

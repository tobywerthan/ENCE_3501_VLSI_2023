*** SPICE deck for cell nand2_1x{sch} from library Lab06
*** Created on Tue Oct 10, 2006 11:35:50
*** Last revised on Sat Nov 11, 2023 19:05:42
*** Written on Sat Nov 11, 2023 19:05:48 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Lab06:nand2_1x{sch}
Mnmos@0 y b net@5 gnd N_50n L=0.6U W=3U
Mnmos@1 net@5 a gnd gnd N_50n L=0.6U W=3U
Mpmos@0 y b vdd vdd P_50n L=0.6U W=6U
Mpmos@1 y a vdd vdd P_50n L=0.6U W=6U
.END

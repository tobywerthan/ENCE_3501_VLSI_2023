*** SPICE deck for cell NOT_gate{lay} from library Werthan_Ring_Oscillator
*** Created on Wed Nov 01, 2023 11:10:59
*** Last revised on Wed Nov 01, 2023 11:19:05
*** Written on Wed Nov 01, 2023 11:19:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NOT_gate{lay}
Mnmos@0 gnd A Y gnd N_1u L=0.6U W=3U AS=7.425P AD=13.5P PS=12.3U PD=23.7U
Mpmos@0 Y A vdd vdd P_1u L=0.6U W=6U AS=18.45P AD=7.425P PS=29.7U PD=12.3U
.END

*** SPICE deck for cell alu{sch} from library Werthan_ALU
*** Created on Sat Nov 11, 2023 11:18:20
*** Last revised on Wed Nov 15, 2023 17:21:56
*** Written on Wed Nov 15, 2023 17:22:02 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_ALU__buftri_c_1x FROM CELL buftri_c_1x{sch}
.SUBCKT Werthan_ALU__buftri_c_1x d en y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@3 net@6 gnd gnd N_1u L=0.6U W=4.2U
Mnmos@1 y en net@3 gnd N_1u L=0.6U W=4.2U
Mnmos@2 net@54 en gnd gnd N_1u L=0.6U W=1.8U
Mnmos@3 net@6 d gnd gnd N_1u L=0.6U W=1.8U
Mpmos@0 net@1 net@54 y vdd P_1u L=0.6U W=6U
Mpmos@1 vdd net@6 net@1 vdd P_1u L=0.6U W=6U
Mpmos@2 vdd en net@54 vdd P_1u L=0.6U W=2.7U
Mpmos@3 vdd d net@6 vdd P_1u L=0.6U W=2.7U
.ENDS Werthan_ALU__buftri_c_1x

*** SUBCIRCUIT Werthan_ALU__fulladder FROM CELL fulladder{sch}
.SUBCKT Werthan_ALU__fulladder a b c cout s
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 a gnd gnd N_1u L=0.6U W=2.4U
Mnmos@1 net@1 b gnd gnd N_1u L=0.6U W=2.4U
Mnmos@2 coutb c net@1 gnd N_1u L=0.6U W=2.4U
Mnmos@3 net@11 a gnd gnd N_1u L=0.6U W=2.4U
Mnmos@4 coutb b net@11 gnd N_1u L=0.6U W=2.4U
Mnmos@5 net@23 a gnd gnd N_1u L=0.6U W=2.4U
Mnmos@6 net@23 b gnd gnd N_1u L=0.6U W=2.4U
Mnmos@7 net@23 c gnd gnd N_1u L=0.6U W=2.4U
Mnmos@8 sb coutb net@23 gnd N_1u L=0.6U W=2.4U
Mnmos@9 net@33 a gnd gnd N_1u L=0.6U W=2.4U
Mnmos@10 net@32 b net@33 gnd N_1u L=0.6U W=2.4U
Mnmos@11 sb c net@32 gnd N_1u L=0.6U W=2.4U
Mnmos@12 cout coutb gnd gnd N_1u L=0.6U W=2.4U
Mnmos@13 s sb gnd gnd N_1u L=0.6U W=2.4U
Mpmos@1 net@92 c sb vdd P_1u L=0.6U W=4.8U
Mpmos@2 net@90 b net@92 vdd P_1u L=0.6U W=4.8U
Mpmos@3 vdd a net@90 vdd P_1u L=0.6U W=4.8U
Mpmos@4 net@94 coutb sb vdd P_1u L=0.6U W=4.8U
Mpmos@5 vdd b net@94 vdd P_1u L=0.6U W=4.8U
Mpmos@6 vdd c net@94 vdd P_1u L=0.6U W=4.8U
Mpmos@7 vdd a net@94 vdd P_1u L=0.6U W=4.8U
Mpmos@8 vdd coutb cout vdd P_1u L=0.6U W=4.8U
Mpmos@9 vdd a net@95 vdd P_1u L=0.6U W=4.8U
Mpmos@10 net@95 b coutb vdd P_1u L=0.6U W=4.8U
Mpmos@11 vdd a net@111 vdd P_1u L=0.6U W=4.8U
Mpmos@12 vdd b net@111 vdd P_1u L=0.6U W=4.8U
Mpmos@13 net@111 c coutb vdd P_1u L=0.6U W=4.8U
Mpmos@14 vdd sb s vdd P_1u L=0.6U W=4.8U
.ENDS Werthan_ALU__fulladder

*** SUBCIRCUIT Werthan_ALU__inv_1x FROM CELL inv_1x{sch}
.SUBCKT Werthan_ALU__inv_1x a y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y a gnd gnd N_1u L=0.6U W=2.1U
Mpmos@0 vdd a y vdd P_1u L=0.6U W=3U
.ENDS Werthan_ALU__inv_1x

*** SUBCIRCUIT Werthan_ALU__mux2_c_1x FROM CELL mux2_c_1x{sch}
.SUBCKT Werthan_ALU__mux2_c_1x d0 d1 s y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@3 d1 gnd gnd N_1u L=0.6U W=1.8U
Mnmos@1 net@4 d0 gnd gnd N_1u L=0.6U W=1.8U
Mnmos@2 net@5 s net@3 gnd N_1u L=0.6U W=1.8U
Mnmos@3 net@5 sb net@4 gnd N_1u L=0.6U W=1.8U
Mnmos@4 y net@5 gnd gnd N_1u L=0.6U W=2.1U
Mnmos@5 sb s gnd gnd N_1u L=0.6U W=1.8U
Mpmos@0 net@15 sb net@5 vdd P_1u L=0.6U W=2.7U
Mpmos@1 vdd d1 net@15 vdd P_1u L=0.6U W=2.7U
Mpmos@2 net@12 s net@5 vdd P_1u L=0.6U W=2.7U
Mpmos@3 vdd d0 net@12 vdd P_1u L=0.6U W=2.7U
Mpmos@4 vdd net@5 y vdd P_1u L=0.6U W=3U
Mpmos@5 vdd s sb vdd P_1u L=0.6U W=2.7U
.ENDS Werthan_ALU__mux2_c_1x

.global gnd vdd

*** TOP LEVEL CELL: alu{sch}
Xbuftri_c@0 net@368 Enable IB[3] Werthan_ALU__buftri_c_1x
Xbuftri_c@1 net@364 Enable IB[2] Werthan_ALU__buftri_c_1x
Xbuftri_c@2 net@359 Enable IB[1] Werthan_ALU__buftri_c_1x
Xbuftri_c@3 net@353 Enable IB[0] Werthan_ALU__buftri_c_1x
Xfulladde@3 B[0] net@78 net@354 net@27 net@353 Werthan_ALU__fulladder
Xfulladde@4 B[1] net@81 net@27 net@8 net@359 Werthan_ALU__fulladder
Xfulladde@5 B[2] net@75 net@8 net@1 net@364 Werthan_ALU__fulladder
Xfulladde@6 B[3] net@70 net@1 carry net@368 Werthan_ALU__fulladder
Xinv_1x@0 A[3] net@311 Werthan_ALU__inv_1x
Xinv_1x@1 A[2] net@313 Werthan_ALU__inv_1x
Xinv_1x@2 A[1] net@318 Werthan_ALU__inv_1x
Xinv_1x@3 A[0] net@320 Werthan_ALU__inv_1x
Xmux2_c_1@0 A[3] net@311 AddSub net@70 Werthan_ALU__mux2_c_1x
Xmux2_c_1@1 A[2] net@313 AddSub net@75 Werthan_ALU__mux2_c_1x
Xmux2_c_1@2 A[1] net@318 AddSub net@81 Werthan_ALU__mux2_c_1x
Xmux2_c_1@3 A[0] net@320 AddSub net@78 Werthan_ALU__mux2_c_1x
Xmux2_c_1@4 vdd gnd AddSub net@354 Werthan_ALU__mux2_c_1x

* Spice Code nodes in cell cell 'alu{sch}'
.include cmosedu_models.txt
.END

*** SPICE deck for cell 5B_R2R_DAC_delay_sim{sch} from library Werthan_5B_R2R_DAC
*** Created on Thu Sep 28, 2023 14:11:05
*** Last revised on Thu Sep 28, 2023 14:17:24
*** Written on Thu Sep 28, 2023 14:17:33 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_R_Divider__R_Divider FROM CELL Werthan_R_Divider:R_Divider{sch}
.SUBCKT Werthan_R_Divider__R_Divider bot in out
Rresnwell@0 net@2 in 10k
Rresnwell@1 out net@2 10k
Rresnwell@2 out bot 10k
.ENDS Werthan_R_Divider__R_Divider

*** SUBCIRCUIT Werthan_5B_R2R_DAC__5B_R2R_DAC FROM CELL 5B_R2R_DAC{sch}
.SUBCKT Werthan_5B_R2R_DAC__5B_R2R_DAC b0 b1 b2 b3 b4 vout
** GLOBAL gnd
Rresnwell@0 net@0 gnd 10k
XR_Divide@0 net@4 b4 vout Werthan_R_Divider__R_Divider
XR_Divide@1 net@3 b3 net@4 Werthan_R_Divider__R_Divider
XR_Divide@2 net@2 b2 net@3 Werthan_R_Divider__R_Divider
XR_Divide@3 net@1 b1 net@2 Werthan_R_Divider__R_Divider
XR_Divide@4 net@0 b0 net@1 Werthan_R_Divider__R_Divider

* Spice Code nodes in cell cell '5B_R2R_DAC{sch}'
*v4 b4 0
*v3 b3 0
*v2 b2 0
*v1 b1 b0
*vin b0 0 DC 5
*.op
.ENDS Werthan_5B_R2R_DAC__5B_R2R_DAC

.global gnd

*** TOP LEVEL CELL: 5B_R2R_DAC_delay_sim{sch}
Ccap@0 gnd vout 10p
X_5B_R2R_D@0 gnd gnd gnd gnd vin vout Werthan_5B_R2R_DAC__5B_R2R_DAC

* Spice Code nodes in cell cell '5B_R2R_DAC_delay_sim{sch}'
vin vin 0 pulse(0v 2v 1u 1f 1f 3u 6u)
.tran 0 2.4u 0 100p
.END

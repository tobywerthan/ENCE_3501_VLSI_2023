*** SPICE deck for cell Vsph_test{sch} from library HW7Q1
*** Created on Sun Nov 05, 2023 17:06:19
*** Last revised on Sun Nov 05, 2023 19:35:55
*** Written on Sun Nov 05, 2023 19:36:01 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Vsph_test{sch}
Mnmos@0 output input net@19 gnd N_50n L=0.6U W=21U
Mnmos@1 net@19 input gnd gnd N_50n L=0.6U W=21U
Mnmos@2 vdd output net@19 gnd N_50n L=0.6U W=9.333U
Mpmos@0 output input net@16 vdd P_50n L=0.6U W=33U
Mpmos@1 net@16 input vdd vdd P_50n L=0.6U W=25.266U
Mpmos@2 gnd output net@16 vdd P_50n L=0.6U W=33U

* Spice Code nodes in cell cell 'Vsph_test{sch}'
.include cmosedu_models.txt
vdd vdd 0 DC 1V
in in 0 SIN(0.5 0.5 50)
.trans 0 40m
.END

*** SPICE deck for cell ring_oscillator_sim{sch} from library Werthan_DC_to_DC
*** Created on Sat Nov 11, 2023 18:36:27
*** Last revised on Sat Nov 11, 2023 19:16:44
*** Written on Sat Nov 11, 2023 19:19:46 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_DC_to_DC__ring_oscillator FROM CELL ring_oscillator{sch}
.SUBCKT Werthan_DC_to_DC__ring_oscillator En osc osc2
** GLOBAL gnd
** GLOBAL vdd
Ccap@0 gnd net@61 10u
Ccap@1 gnd net@67 10u
Ccap@2 gnd net@73 10u
Mnmos@0 net@61 En net@77 gnd N_50n L=0.6U W=3U
Mnmos@1 net@77 osc gnd gnd N_50n L=0.6U W=3U
Mnmos@2 net@73 net@61 gnd gnd N_50n L=0.6U W=3U
Mnmos@3 net@67 net@73 gnd gnd N_50n L=0.6U W=3U
Mnmos@4 osc2 net@67 gnd gnd N_50n L=0.6U W=3U
Mnmos@5 osc osc2 gnd gnd N_50n L=0.6U W=3U
Mpmos@0 net@61 En vdd vdd P_50n L=0.6U W=6U
Mpmos@1 net@61 osc vdd vdd P_50n L=0.6U W=6U
Mpmos@2 net@73 net@61 vdd vdd P_50n L=0.6U W=6U
Mpmos@3 net@67 net@73 vdd vdd P_50n L=0.6U W=6U
Mpmos@4 osc2 net@67 vdd vdd P_50n L=0.6U W=6U
Mpmos@5 osc osc2 vdd vdd P_50n L=0.6U W=6U
.ENDS Werthan_DC_to_DC__ring_oscillator

.global gnd vdd

*** TOP LEVEL CELL: ring_oscillator_sim{sch}
Xring_osc@0 en osc osc2 Werthan_DC_to_DC__ring_oscillator

* Spice Code nodes in cell cell 'ring_oscillator_sim{sch}'
vdd vdd 0 DC 1v
ven en 0 dc 1v
.tran 0 10
.include cmosedu_models.txt
.END

*** SPICE deck for cell 5B_R2R_DAC_sim{sch} from library Werthan_5B_R2R_DAC
*** Created on Sun Sep 24, 2023 14:59:49
*** Last revised on Tue Sep 26, 2023 16:44:37
*** Written on Tue Sep 26, 2023 16:44:44 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Werthan_5B_R2R_DAC__R_Divider FROM CELL Werthan_5B_R2R_DAC:R_Divider{sch}
.SUBCKT Werthan_5B_R2R_DAC__R_Divider bot in out
Rresnwell@0 net@2 in 10k
Rresnwell@1 out net@2 10k
Rresnwell@2 out bot 10k
.ENDS Werthan_5B_R2R_DAC__R_Divider

*** SUBCIRCUIT Werthan_5B_R2R_DAC__5B_R2R_DAC FROM CELL Werthan_5B_R2R_DAC:5B_R2R_DAC{sch}
.SUBCKT Werthan_5B_R2R_DAC__5B_R2R_DAC b0 b1 b2 b3 b4 vout
** GLOBAL gnd
Rresnwell@0 net@0 gnd 10k
XR_Divide@0 net@4 b4 vout Werthan_5B_R2R_DAC__R_Divider
XR_Divide@1 net@3 b3 net@4 Werthan_5B_R2R_DAC__R_Divider
XR_Divide@2 net@2 b2 net@3 Werthan_5B_R2R_DAC__R_Divider
XR_Divide@3 net@1 b1 net@2 Werthan_5B_R2R_DAC__R_Divider
XR_Divide@4 net@0 b0 net@1 Werthan_5B_R2R_DAC__R_Divider
.ENDS Werthan_5B_R2R_DAC__5B_R2R_DAC

.global gnd

*** TOP LEVEL CELL: Werthan_5B_R2R_DAC:5B_R2R_DAC_sim{sch}
X_5B_R2R_D@0 vin vin gnd gnd gnd vout Werthan_5B_R2R_DAC__5B_R2R_DAC
.END
